user@machine.23855:1689094962