user@machine.15452:1691585023